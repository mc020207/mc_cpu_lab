`ifndef __CORE_SV
`define __CORE_SV
`ifdef VERILATOR
`include "include/common.sv"
`include "include/pipes.sv"
`include "pipeline/regfile/regfile.sv"
`include "pipeline/fetch/fetch.sv"
`include "pipeline/decode/decode.sv"
`include "pipeline/execute/execute.sv"
`include "pipeline/memory/memory.sv"
`include "pipeline/regfile/csr.sv"
`else

`endif

module core 
	import common::*;
	import pipes::*;(
	input logic clk, reset,
	output ibus_req_t  ireq,
	input  ibus_resp_t iresp,
	output dbus_req_t  dreq,
	input  dbus_resp_t dresp,
	input logic trint, swint, exint
);
	fetch_data_t dataF;
	decode_data_t dataD;
	excute_data_t dataE;
	memory_data_t dataM;
	creg_addr_t ra1,ra2;
	word_t rd1,rd2;
	u1 stopf,stopd,stope,stopm,branch;
	u1 flushde,flushall;
	u64 jump;
	tran_t trane,tranm,tranw;
	u12 csrra;
	word_t csrrd;
	u64 csrpc;
	fetch fetch(
		.clk,.reset,
		.ireq,.iresp,
		.branch,.jump,
		.stopd,.stope,.stopm,
		.dataF,.stopf,.flushde,.flushall,.csrpc
	);
	decode decode (
		.clk,.reset,
		.dataF,.dataD,
		.ra1,.ra2,.rd1,.rd2,
		.branch,
		.trane,.tranm,.tranw,
		.stopd,.stope,.stopm,
		.csrra,.csrrd,.flushde
	);
	regfile regfile(
		.clk, .reset,
		.ra1,.ra2,.rd1,.rd2,
		.wvalid(dataM.ctl.regwrite&&dataM.valid),
		.wa(dataM.dst),
		.wd(dataM.result)
	);
	csr csrreg(
		.clk,.reset,
		.ra(csrra),.rd(csrrd),
		.dataM,.csrpc,.trint,.swint,.exint,
		.stopf,.stopm,.flushde,.flushall
	);
	execute execute(
		.clk,.reset,
		.dataD,.dataE,
		.branch,.jump,
		.trane,.stope,.stopm,.flushde
	);
	memory memory(
		.clk,.reset,
		.dataE,.dataM(dataM),
		.dreq,.dresp,
		.tranm,.stopm,.flushde,.flushall
	);
	logic skip;
	assign skip=(dataM.ctl.op==SD||dataM.ctl.op==LD)&&dataM.addr[31]==0;
	assign tranw.dst=(dataM.ctl.regwrite&dataM.valid&&(dataM.error==0))?dataM.dst:0;
	assign tranw.data=dataM.result;
	assign tranw.ismem=1;
`ifdef VERILATOR
	DifftestInstrCommit DifftestInstrCommit(
		.clock              (clk),
		.coreid             (0),
		.index              (0),
		.valid              (~reset&&dataM.valid&&(dataM.error==0)),
		.pc                 (dataM.pc),
		.instr              (dataM.raw_instr),
		.skip               (skip),
		.isRVC              (0),
		.scFailed           (0),
		.wen                (dataM.ctl.regwrite),
		.wdest              ({3'b0,dataM.dst}),
		.wdata              (dataM.result)
	);
	      
	DifftestArchIntRegState DifftestArchIntRegState (
		.clock              (clk),
		.coreid             (0),
		.gpr_0              (regfile.regs_nxt[0]),
		.gpr_1              (regfile.regs_nxt[1]),
		.gpr_2              (regfile.regs_nxt[2]),
		.gpr_3              (regfile.regs_nxt[3]),
		.gpr_4              (regfile.regs_nxt[4]),
		.gpr_5              (regfile.regs_nxt[5]),
		.gpr_6              (regfile.regs_nxt[6]),
		.gpr_7              (regfile.regs_nxt[7]),
		.gpr_8              (regfile.regs_nxt[8]),
		.gpr_9              (regfile.regs_nxt[9]),
		.gpr_10             (regfile.regs_nxt[10]),
		.gpr_11             (regfile.regs_nxt[11]),
		.gpr_12             (regfile.regs_nxt[12]),
		.gpr_13             (regfile.regs_nxt[13]),
		.gpr_14             (regfile.regs_nxt[14]),
		.gpr_15             (regfile.regs_nxt[15]),
		.gpr_16             (regfile.regs_nxt[16]),
		.gpr_17             (regfile.regs_nxt[17]),
		.gpr_18             (regfile.regs_nxt[18]),
		.gpr_19             (regfile.regs_nxt[19]),
		.gpr_20             (regfile.regs_nxt[20]),
		.gpr_21             (regfile.regs_nxt[21]),
		.gpr_22             (regfile.regs_nxt[22]),
		.gpr_23             (regfile.regs_nxt[23]),
		.gpr_24             (regfile.regs_nxt[24]),
		.gpr_25             (regfile.regs_nxt[25]),
		.gpr_26             (regfile.regs_nxt[26]),
		.gpr_27             (regfile.regs_nxt[27]),
		.gpr_28             (regfile.regs_nxt[28]),
		.gpr_29             (regfile.regs_nxt[29]),
		.gpr_30             (regfile.regs_nxt[30]),
		.gpr_31             (regfile.regs_nxt[31])
	);
	      
	DifftestTrapEvent DifftestTrapEvent(
		.clock              (clk),
		.coreid             (0),
		.valid              (0),
		.code               (0),
		.pc                 (0),
		.cycleCnt           (0),
		.instrCnt           (0)
	);
	      
	DifftestCSRState DifftestCSRState(
		.clock              (clk),
		.coreid             (0),
		.priviledgeMode     (csrreg.mode_nxt),
		.mstatus            (csrreg.regs_nxt.mstatus),
		.sstatus            (csrreg.regs_nxt.mstatus & 64'h800000030001e000),
		.mepc               (csrreg.regs_nxt.mepc),
		.sepc               (0),
		.mtval              (csrreg.regs_nxt.mtval),
		.stval              (0),
		.mtvec              (csrreg.regs_nxt.mtvec),
		.stvec              (0),
		.mcause             (csrreg.regs_nxt.mcause),
		.scause             (0),
		.satp               (0),
		.mip                (csrreg.regs_nxt.mip),
		.mie                (csrreg.regs_nxt.mie),
		.mscratch           (csrreg.regs_nxt.mscratch),
		.sscratch           (0),
		.mideleg            (0),
		.medeleg            (0)
	);
	      
	DifftestArchFpRegState DifftestArchFpRegState(
		.clock              (clk),
		.coreid             (0),
		.fpr_0              (0),
		.fpr_1              (0),
		.fpr_2              (0),
		.fpr_3              (0),
		.fpr_4              (0),
		.fpr_5              (0),
		.fpr_6              (0),
		.fpr_7              (0),
		.fpr_8              (0),
		.fpr_9              (0),
		.fpr_10             (0),
		.fpr_11             (0),
		.fpr_12             (0),
		.fpr_13             (0),
		.fpr_14             (0),
		.fpr_15             (0),
		.fpr_16             (0),
		.fpr_17             (0),
		.fpr_18             (0),
		.fpr_19             (0),
		.fpr_20             (0),
		.fpr_21             (0),
		.fpr_22             (0),
		.fpr_23             (0),
		.fpr_24             (0),
		.fpr_25             (0),
		.fpr_26             (0),
		.fpr_27             (0),
		.fpr_28             (0),
		.fpr_29             (0),
		.fpr_30             (0),
		.fpr_31             (0)
	);
	
`endif
endmodule
`endif